RAM_OUTENAB_MUX_inst : RAM_OUTENAB_MUX PORT MAP (
		data0	 => data0_sig,
		data1	 => data1_sig,
		sel	 => sel_sig,
		result	 => result_sig
	);
