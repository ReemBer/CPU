INCS_LOAD_BUSTRI_inst : INCS_LOAD_BUSTRI PORT MAP (
		data	 => data_sig,
		enabledt	 => enabledt_sig,
		tridata	 => tridata_sig
	);
