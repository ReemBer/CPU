STACK_POINTER_ASYNC_SET_COMPARATOR_inst : STACK_POINTER_ASYNC_SET_COMPARATOR PORT MAP (
		dataa	 => dataa_sig,
		AeB	 => AeB_sig
	);
