INDIRECT_ADDRESSING_MUX_inst : INDIRECT_ADDRESSING_MUX PORT MAP (
		data0x	 => data0x_sig,
		data1x	 => data1x_sig,
		sel	 => sel_sig,
		result	 => result_sig
	);
