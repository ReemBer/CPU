IP_REGISTER_inst : IP_REGISTER PORT MAP (
		clock	 => clock_sig,
		data	 => data_sig,
		q	 => q_sig
	);
