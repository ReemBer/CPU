ALU_RESULT_BUSTRI_inst : ALU_RESULT_BUSTRI PORT MAP (
		data	 => data_sig,
		enabledt	 => enabledt_sig,
		tridata	 => tridata_sig
	);
