STACK_POINTER_DECODER_inst : STACK_POINTER_DECODER PORT MAP (
		data	 => data_sig,
		eq0	 => eq0_sig,
		eq1	 => eq1_sig,
		eq2	 => eq2_sig,
		eq3	 => eq3_sig,
		eq4	 => eq4_sig
	);
