SRA_DISTANCE_REGISTER_inst : SRA_DISTANCE_REGISTER PORT MAP (
		clock	 => clock_sig,
		data	 => data_sig,
		enable	 => enable_sig,
		q	 => q_sig
	);
