RW_RAM_BUSTRI_inst : RW_RAM_BUSTRI PORT MAP (
		data	 => data_sig,
		enabledt	 => enabledt_sig,
		enabletr	 => enabletr_sig,
		result	 => result_sig,
		tridata	 => tridata_sig
	);
