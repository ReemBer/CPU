ALU_NOTZ_REGISTER_inst : ALU_NOTZ_REGISTER PORT MAP (
		clock	 => clock_sig,
		data	 => data_sig,
		enable	 => enable_sig,
		q	 => q_sig
	);
