ALU_NOTZ_OUT_MUX_inst : ALU_NOTZ_OUT_MUX PORT MAP (
		data0x	 => data0x_sig,
		data1x	 => data1x_sig,
		sel	 => sel_sig,
		result	 => result_sig
	);
