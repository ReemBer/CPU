CPU_CYCLE_COUNTER_inst : CPU_CYCLE_COUNTER PORT MAP (
		aclr	 => aclr_sig,
		clk_en	 => clk_en_sig,
		clock	 => clock_sig,
		sclr	 => sclr_sig,
		q	 => q_sig
	);
