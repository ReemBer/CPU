RAM_ADDRESS_BUSTRI_inst : RAM_ADDRESS_BUSTRI PORT MAP (
		data	 => data_sig,
		enabledt	 => enabledt_sig,
		tridata	 => tridata_sig
	);
