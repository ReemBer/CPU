NEW_IP_TEST_inst : NEW_IP_TEST PORT MAP (
		clk_en	 => clk_en_sig,
		clock	 => clock_sig,
		data	 => data_sig,
		sload	 => sload_sig,
		q	 => q_sig
	);
