ALU_SRA_SHIFT_REGISTER_inst : ALU_SRA_SHIFT_REGISTER PORT MAP (
		data	 => data_sig,
		distance	 => distance_sig,
		result	 => result_sig,
		underflow	 => underflow_sig
	);
