Z_FLAG_OR_inst : Z_FLAG_OR PORT MAP (
		data	 => data_sig,
		result	 => result_sig
	);
