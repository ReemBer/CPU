ALU_INPUT_BUSTRI_inst : ALU_INPUT_BUSTRI PORT MAP (
		data	 => data_sig,
		enabledt	 => enabledt_sig,
		tridata	 => tridata_sig
	);
