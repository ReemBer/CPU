RAM_DIRECT_ADDRESS_inst : RAM_DIRECT_ADDRESS PORT MAP (
		clock	 => clock_sig,
		data	 => data_sig,
		enable	 => enable_sig,
		q	 => q_sig
	);
