STACK_POINTER_COUNTER_inst : STACK_POINTER_COUNTER PORT MAP (
		aclr	 => aclr_sig,
		aset	 => aset_sig,
		clock	 => clock_sig,
		updown	 => updown_sig,
		q	 => q_sig
	);
