STACK_OUT_BUSTRI_inst : STACK_OUT_BUSTRI PORT MAP (
		data	 => data_sig,
		enabledt	 => enabledt_sig,
		tridata	 => tridata_sig
	);
