GENERAL_REGISTER_READ_BUSTRI_inst : GENERAL_REGISTER_READ_BUSTRI PORT MAP (
		data	 => data_sig,
		enabledt	 => enabledt_sig,
		tridata	 => tridata_sig
	);
