CPU_DATA_BUS_OUT_MUX_inst : CPU_DATA_BUS_OUT_MUX PORT MAP (
		data0x	 => data0x_sig,
		data1x	 => data1x_sig,
		sel	 => sel_sig,
		result	 => result_sig
	);
