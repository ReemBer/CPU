C_FLAG_inst : C_FLAG PORT MAP (
		aclr	 => aclr_sig,
		aset	 => aset_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
