ALU_SRA_REGISTER_inst : ALU_SRA_REGISTER PORT MAP (
		clock	 => clock_sig,
		data	 => data_sig,
		enable	 => enable_sig,
		q	 => q_sig
	);
