IP_COUNTER_inst : IP_COUNTER PORT MAP (
		clock	 => clock_sig,
		data	 => data_sig,
		sload	 => sload_sig,
		q	 => q_sig
	);
