NOTZ_XOR_inst : NOTZ_XOR PORT MAP (
		data	 => data_sig,
		result	 => result_sig
	);
