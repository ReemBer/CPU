CPU_CYCLE_COUNTER_inst : CPU_CYCLE_COUNTER PORT MAP (
		clock	 => clock_sig,
		sclr	 => sclr_sig,
		q	 => q_sig
	);
