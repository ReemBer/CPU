ALU_OUTPUT_BUSTRI_inst : ALU_OUTPUT_BUSTRI PORT MAP (
		data	 => data_sig,
		enabledt	 => enabledt_sig,
		tridata	 => tridata_sig
	);
