ALU_NXOR_FIRST_REGISTER_inst : ALU_NXOR_FIRST_REGISTER PORT MAP (
		clock	 => clock_sig,
		data	 => data_sig,
		enable	 => enable_sig,
		q	 => q_sig
	);
