NXOR_INVERTOR_inst : NXOR_INVERTOR PORT MAP (
		data	 => data_sig,
		result	 => result_sig
	);
