lpm_ff0_inst : lpm_ff0 PORT MAP (
		aclr	 => aclr_sig,
		aset	 => aset_sig,
		clock	 => clock_sig,
		data	 => data_sig,
		q	 => q_sig
	);
