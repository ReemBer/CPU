STACK_POINTER_ASYNC_CLEAR_COMPARATOR_inst : STACK_POINTER_ASYNC_CLEAR_COMPARATOR PORT MAP (
		dataa	 => dataa_sig,
		AeB	 => AeB_sig
	);
