STACK_REGISTER_inst : STACK_REGISTER PORT MAP (
		clock	 => clock_sig,
		data	 => data_sig,
		enable	 => enable_sig,
		q	 => q_sig
	);
