COMMAND_WORD_BUFFER_inst : COMMAND_WORD_BUFFER PORT MAP (
		clock	 => clock_sig,
		data	 => data_sig,
		q	 => q_sig
	);
