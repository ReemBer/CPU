IP_inst : IP PORT MAP (
		clk_en	 => clk_en_sig,
		clock	 => clock_sig,
		data	 => data_sig,
		sload	 => sload_sig,
		q	 => q_sig
	);
