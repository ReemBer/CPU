NOTZ_INVERTOR_inst : NOTZ_INVERTOR PORT MAP (
		data	 => data_sig,
		result	 => result_sig
	);
