IP_TEST_ENTITY_inst : IP_TEST_ENTITY PORT MAP (
		clock	 => clock_sig,
		data	 => data_sig,
		sload	 => sload_sig,
		q	 => q_sig
	);
