NXOR_SECOND_OPERAND_ID_MUX_inst : NXOR_SECOND_OPERAND_ID_MUX PORT MAP (
		data0x	 => data0x_sig,
		data1x	 => data1x_sig,
		sel	 => sel_sig,
		result	 => result_sig
	);
