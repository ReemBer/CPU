IP_BUSTRI_inst : IP_BUSTRI PORT MAP (
		data	 => data_sig,
		enabledt	 => enabledt_sig,
		tridata	 => tridata_sig
	);
