IP_REG_TEST_inst : IP_REG_TEST PORT MAP (
		clock	 => clock_sig,
		data	 => data_sig,
		q	 => q_sig
	);
